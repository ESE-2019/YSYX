// module bpu
//   import OoO_pkg::*;
// (
//     input logic clock,
//     input logic reset,

//     input logic [31:0] pc
// );

// endmodule
