`default_nettype none

module ysyx_24080006_pc
  import OoO_pkg::*;
(
    input logic clock,
    input logic reset
);


endmodule

`default_nettype wire
