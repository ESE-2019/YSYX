// module bpu
//   import ysyx_24080006_pkg::*;
// (
//     input logic clock,
//     input logic reset,

//     input logic [31:0] pc
// );

// endmodule
